LIBRARY ieee;
USE ieee.std_logic_1164.all;


PACKAGE aux_package IS

	COMPONENT top IS
	GENERIC (n : INTEGER);
	PORT (  cin : IN STD_LOGIC;
			sel : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
			X,Y: IN STD_LOGIC_VECTOR (n-1 DOWNTO 0);
		    result: OUT STD_LOGIC_VECTOR(n downto 0));
	END COMPONENT;

	COMPONENT FA IS
	PORT (  xi,yi,cin : IN STD_LOGIC;
			s,cout: OUT STD_LOGIC);
	END COMPONENT;

	COMPONENT selector IS
	GENERIC (n : INTEGER := 8);
	PORT (     in1:  IN STD_LOGIC_VECTOR(n DOWNTO 0);
			  in2: IN STD_LOGIC_VECTOR(8 DOWNTO 0);
		     sel: IN STD_LOGIC_VECTOR(1 downto 0);
             output: OUT STD_LOGIC_VECTOR(n DOWNTO 0));
	END COMPONENT;
	
	COMPONENT Barrel IS
	PORT (  x: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			y: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
			output: OUT STD_LOGIC_VECTOR(8 downto 0));
	END COMPONENT;
	
	COMPONENT MuxCombined IS
	GENERIC (n : INTEGER);
	PORT (  x1,x2: IN STD_LOGIC_VECTOR (n-1 DOWNTO 0);
			sel: IN STD_LOGIC;
			output: OUT STD_LOGIC_VECTOR(n-1 downto 0));
	END COMPONENT;
	
	COMPONENT mux2on1 IS
	PORT (  in1,in2,sel: IN STD_LOGIC;
			output: OUT STD_LOGIC);
	END COMPONENT;
	
	
	COMPONENT AdderTwo IS
	GENERIC (n : INTEGER);
	PORT (   cin: IN STD_LOGIC;
			 x,y: IN STD_LOGIC_VECTOR (n-1 DOWNTO 0);
			 sel : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
             s: OUT STD_LOGIC_VECTOR(n DOWNTO 0));
	END COMPONENT;
  
END aux_package;

