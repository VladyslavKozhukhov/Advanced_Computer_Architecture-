 LIBRARY IEEE;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;
USE ieee.std_logic_unsigned.all;
USE work.aux_package_cond.all;

ENTITY cond_tb IS
	CONSTANT n : INTEGER := 8;
END cond_tb;
 
 
architecture cond_Testbench OF cond_tb IS
SIGNAL rst,ena,clk: STD_LOGIC;
	SIGNAL din: STD_LOGIC_VECTOR (n-1 DOWNTO 0);
	SIGNAL condd: INTEGER range 0 to 3;
	SIGNAL	detector : std_logic;
	SIGNAL	D_prev :  std_logic_vector(n-1 downto 0);
BEGIN

	L0 : Cond PORT MAP(rst,ena,clk,D_prev,condd,din,detector);
tb_ena : process
			begin
			ena<='0';
			wait for 20 us;

			ena<='1';
			
			wait;
        end process tb_ena;
		
	tb_cond : process
		begin
				condd<=0;		

			wait;
			
	end process tb_cond;

        tb_clk : process
			begin 
			clk<='0';
			wait for 5 us;
			clk<='1';
			wait for 5 us;
        end process tb_clk;
		
		tb_rst : process
			begin 
			rst<='1';
			wait for 10 us;
			rst<='0';
			wait;
        end process tb_rst;
		
		
    tb_din : process
		begin
			D_prev <= "00000000";
			din<="00000001";
			wait for 10 us;
			D_prev <= "00000001";
			din<="00000010";

			wait for 10 us;
			D_prev <= "00000010";
			din<="00000011";

			wait for 10 us;
			din <= "00000011"; 
			D_prev<="00000011";
			wait for 10 us;
			D_prev <= "00000100";
			din<="00000101";
			
			wait ;
        end process tb_din;
		

  
  
END cond_Testbench;