LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
---finish  sll srl 
ENTITY MIPS IS

	PORT( reset, clock					: IN 	STD_LOGIC;
	-----------------------------------------------------------
		IsTEST: OUT std_logic;
		sw_8_run: IN std_logic; -- for IO
		sw_0_7 : IN std_logic_vector(7 DOWNTO 0); --for IO
		HI_OUT: OUT std_logic_vector(7 DOWNTO 0); -- for IO
		LO_OUT: OUT std_logic_vector(7 DOWNTO 0); -- for IO
		SEG0_OUT, SEG1_OUT: OUT std_logic_vector(6 DOWNTO 0); -- for IO
		SEG2_OUT, SEG3_OUT: OUT std_logic_vector(6 DOWNTO 0); -- for IO
		PORT_LEDG: OUT std_logic_vector(7 DOWNTO 0);-- for IO
		PORT_LEDR: OUT std_logic_vector(7 DOWNTO 0);-- for IO

	-----------------------------------------------------------
		-- Output important signals to pins for easy display in Simulator
		PC								: OUT  STD_LOGIC_VECTOR( 9 DOWNTO 0 );
		ALU_result_out, read_data_1_out, read_data_2_out, write_data_out,	
     	Instruction_out					: OUT 	STD_LOGIC_VECTOR( 31 DOWNTO 0 );
		Branch_out, Zero_out, Memwrite_out, 
		Regwrite_out					: OUT 	STD_LOGIC );
END 	MIPS;

ARCHITECTURE structure OF MIPS IS

	COMPONENT Ifetch
   	     PORT(	Instruction			: OUT 	STD_LOGIC_VECTOR( 31 DOWNTO 0 );
        		PC_plus_4_out 		: OUT  	STD_LOGIC_VECTOR( 9 DOWNTO 0 );
				bubble_out			: OUT	STD_LOGIC;----
				IsSpecialAddr		: IN    std_logic;
        		Add_result 			: IN 	STD_LOGIC_VECTOR( 7 DOWNTO 0 );
        		Branch 				: IN 	STD_LOGIC;
        		Zero 				: IN 	STD_LOGIC;
        		Jump 				: IN 	STD_LOGIC;
				sw_8_run			: IN 	std_logic;
        		PC_out 				: OUT 	STD_LOGIC_VECTOR( 9 DOWNTO 0 );
        		clock,reset 		: IN 	STD_LOGIC );
	END COMPONENT; 

	COMPONENT Idecode
 	     PORT(	read_data_1 		: OUT 	STD_LOGIC_VECTOR( 31 DOWNTO 0 );
        		read_data_2 		: OUT 	STD_LOGIC_VECTOR( 31 DOWNTO 0 );
        		Instruction 		: IN 	STD_LOGIC_VECTOR( 31 DOWNTO 0 );
        		read_data 			: IN 	STD_LOGIC_VECTOR( 31 DOWNTO 0 );
        		ALU_result 			: IN 	STD_LOGIC_VECTOR( 31 DOWNTO 0 );
        		RegWrite, MemtoReg 	: IN 	STD_LOGIC;
        		RegDst 				: IN 	STD_LOGIC;
				bubble_out			: IN  	STD_LOGIC;---
        		Sign_extend 		: OUT 	STD_LOGIC_VECTOR( 31 DOWNTO 0 );
				IsSpecialAddr		: OUT    std_logic;
				IsTEST: OUT std_logic;
				addrOfIO    :OUT STD_LOGIC_VECTOR(11 downto 0);--addr of IO
        		clock, reset		: IN 	STD_LOGIC );
	END COMPONENT;

	COMPONENT control
	     PORT( 	Opcode 				: IN 	STD_LOGIC_VECTOR( 5 DOWNTO 0 );
             	RegDst 				: OUT 	STD_LOGIC;
             	ALUSrc 				: OUT 	STD_LOGIC;
             	MemtoReg 			: OUT 	STD_LOGIC;
             	RegWrite 			: OUT 	STD_LOGIC;
             	MemRead 			: OUT 	STD_LOGIC;
             	MemWrite 			: OUT 	STD_LOGIC;
             	Branch 				: OUT 	STD_LOGIC;
             	ALUop 				: OUT 	STD_LOGIC_VECTOR( 1 DOWNTO 0 );
				Jump				: OUT 	STD_LOGIC; 
				ICommand	: OUT 	STD_LOGIC_VECTOR( 3 DOWNTO 0 );
	SLWCommand	: OUT 	STD_LOGIC_VECTOR( 3 DOWNTO 0 );
	IsICommand  : OUT 	STD_LOGIC;
	IsSWCommand  : OUT 	STD_LOGIC;
             	clock, reset		: IN 	STD_LOGIC );
	END COMPONENT;

	COMPONENT  Execute
   	     PORT(	Read_data_1 		: IN 	STD_LOGIC_VECTOR( 31 DOWNTO 0 );
                Read_data_2 		: IN 	STD_LOGIC_VECTOR( 31 DOWNTO 0 );
               	Sign_Extend 		: IN 	STD_LOGIC_VECTOR( 31 DOWNTO 0 );
               	Function_opcode		: IN 	STD_LOGIC_VECTOR( 5 DOWNTO 0 );
               	ALUOp 				: IN 	STD_LOGIC_VECTOR( 1 DOWNTO 0 );
               	ALUSrc 				: IN 	STD_LOGIC;
               	Zero 				: OUT	STD_LOGIC;
               	ALU_Result 			: OUT	STD_LOGIC_VECTOR( 31 DOWNTO 0 );
               	Add_Result 			: OUT	STD_LOGIC_VECTOR( 7 DOWNTO 0 );
               	PC_plus_4 			: IN 	STD_LOGIC_VECTOR( 9 DOWNTO 0 );
				ICommand	: IN 	STD_LOGIC_VECTOR( 3 DOWNTO 0 );
	SLWCommand	: IN 	STD_LOGIC_VECTOR( 3 DOWNTO 0 );
	IsICommand  : IN 	STD_LOGIC;
	IsSWCommand  : IN 	STD_LOGIC;
				shiftValue			: IN    STD_LOGIC_VECTOR( 4 DOWNTO 0 );
               	clock, reset		: IN 	STD_LOGIC );
	END COMPONENT;


	COMPONENT dmemory
	     PORT(	read_data 			: OUT 	STD_LOGIC_VECTOR( 31 DOWNTO 0 );
        		address 			: IN 	STD_LOGIC_VECTOR( 9 DOWNTO 0 );
        		write_data 			: IN 	STD_LOGIC_VECTOR( 31 DOWNTO 0 );
        		MemRead, Memwrite 	: IN 	STD_LOGIC;
				SpecialAddr         : IN 	STD_LOGIC;
				SpecialData         : IN    std_logic_vector(7 DOWNTO 0);
				IsSpecialAddr		: IN    std_logic;
				Seven_Seg			: OUT 	STD_LOGIC_VECTOR( 15 downto 0 );
				PORT_LEDG: OUT std_logic_vector(7 DOWNTO 0);-- for IO
				PORT_LEDR: OUT std_logic_vector(7 DOWNTO 0);-- for IO
				addrOfIO    :IN STD_LOGIC_VECTOR(11 downto 0);--addr of IO

        		Clock,reset			: IN 	STD_LOGIC );
	END COMPONENT;
		-----------------------------------------------------------------
COMPONENT sevenSegment IS
	PORT (
		HI, LO : IN std_logic_vector(7 DOWNTO 0);
		----------------------------------------
		SEG0_OUT, SEG1_OUT: OUT std_logic_vector(6 DOWNTO 0);
		SEG2_OUT, SEG3_OUT: OUT std_logic_vector(6 DOWNTO 0)
	);
END COMPONENT;

COMPONENT BCD 
	port ( 	Binary: 	in  std_logic_vector(3 downto 0);
			En:			in  std_logic;
			Hex_out:	out std_logic_vector(6 downto 0));
end COMPONENT;
	
COMPONENT Ndff
	 GENERIC ( N: integer := 8);
	 PORT (	d					: in std_logic_vector(N-1 downto 0);
			clk					: in std_logic;
			rst					: in std_logic;
			q					: out std_logic_vector(N-1 downto 0) );
END COMPONENT;
--------------------------------------
					-- declare signals used to connect VHDL components
	SIGNAL PC_plus_4 		: STD_LOGIC_VECTOR( 9 DOWNTO 0 );
	SIGNAL read_data_1 		: STD_LOGIC_VECTOR( 31 DOWNTO 0 );
	SIGNAL read_data_2 		: STD_LOGIC_VECTOR( 31 DOWNTO 0 );
	SIGNAL Sign_Extend 		: STD_LOGIC_VECTOR( 31 DOWNTO 0 );
	SIGNAL Add_result 		: STD_LOGIC_VECTOR( 7 DOWNTO 0 );
	SIGNAL ALU_result 		: STD_LOGIC_VECTOR( 31 DOWNTO 0 );
	SIGNAL read_data 		: STD_LOGIC_VECTOR( 31 DOWNTO 0 );
	SIGNAL ALUSrc 			: STD_LOGIC;
	SIGNAL Branch 			: STD_LOGIC;
	SIGNAL Jump				: STD_LOGIC;
	SIGNAL SpecialAddr      : STD_LOGIC;
	SIGNAL IsSpecialAddr    : STD_LOGIC;
	SIGNAL ICommand	        : STD_LOGIC_VECTOR( 3 DOWNTO 0 );
	SIGNAL shiftValue		: STD_LOGIC_VECTOR( 4 DOWNTO 0 );
	SIGNAL IsICommand       : STD_LOGIC;
	SIGNAL	SLWCommand	:  	STD_LOGIC_VECTOR( 3 DOWNTO 0 );

	SIGNAL IsSWCommand: STD_LOGIC;
	SIGNAL RegDst 			: STD_LOGIC;
	SIGNAL Regwrite 		: STD_LOGIC;
	SIGNAL Zero 			: STD_LOGIC;
	SIGNAL MemWrite 		: STD_LOGIC;
	SIGNAL MemtoReg 		: STD_LOGIC;
	SIGNAL MemRead 			: STD_LOGIC;
	SIGNAL ALUop 			: STD_LOGIC_VECTOR(  1 DOWNTO 0 );
	SIGNAL Instruction		: STD_LOGIC_VECTOR( 31 DOWNTO 0 );
	SIGNAL 			addrOfIO    : STD_LOGIC_VECTOR(11 downto 0);--addr of IO
	SIGNAL address_tmp 			:STD_LOGIC_VECTOR( 9 DOWNTO 0 );

		--seven seg vars--------
	SIGNAL ssg0_out					: STD_LOGIC_VECTOR( 6 DOWNTO 0 );
	SIGNAL ssg1_out					: STD_LOGIC_VECTOR( 6 DOWNTO 0 );
	SIGNAL ssg2_out					: STD_LOGIC_VECTOR( 6 DOWNTO 0 );
	SIGNAL ssg3_out					: STD_LOGIC_VECTOR( 6 DOWNTO 0 );
	SIGNAL Seven_Seg				: STD_LOGIC_VECTOR( 15 DOWNTO 0 );
	signal seg_signal_0 : STD_LOGIC_VECTOR( 6 DOWNTO 0 );
	signal seg_signal_1 : STD_LOGIC_VECTOR( 6 DOWNTO 0 );
	signal seg_signal_2 : STD_LOGIC_VECTOR( 6 DOWNTO 0 );
	signal seg_signal_3 : STD_LOGIC_VECTOR( 6 DOWNTO 0 );
	signal the_one						: STD_LOGIC;
   -------------------------------------
	SIGNAL bubble_delay			: STD_LOGIC_VECTOR	(0 downto 0);

BEGIN
					-- copy important signals to output pins for easy 
					-- display in Simulator
   Instruction_out 	<= Instruction;
   ALU_result_out 	<= ALU_result;
   read_data_1_out 	<= read_data_1;
   read_data_2_out 	<= read_data_2;
   write_data_out  	<= read_data WHEN MemtoReg = '1' ELSE ALU_result;
   Branch_out 		<= Branch;
   Zero_out 		<= Zero;
   RegWrite_out 	<= RegWrite;
   MemWrite_out 	<= MemWrite;	
   -------------------------------------
   the_one <= '1';
   SEG0_OUT <= ssg0_out;--seg_signal_0;
   SEG1_OUT <=ssg1_out;-- seg_signal_1;
   SEG2_OUT <= ssg2_out;--seg_signal_2;
   SEG3_OUT <=ssg3_out;-- seg_signal_3;
   
   
   address_tmp<= ALU_Result (9 DOWNTO 2)&"00";
   
   
   ---------------------------------------
					-- connect the 5 MIPS components   
  IFE : Ifetch
	PORT MAP (	Instruction 	=> Instruction,
    	    	PC_plus_4_out 	=> PC_plus_4,
				bubble_out		=> bubble_delay(0),---
				IsSpecialAddr   =>IsSpecialAddr,---
				Add_result 		=> Add_result,
				Branch 			=> Branch,
				Zero 			=> Zero,
				Jump 			=> Jump, 
				sw_8_run	    => sw_8_run,
				PC_out 			=> PC,        		
				clock 			=> clock,  
				reset 			=> reset );

   ID : Idecode
   	PORT MAP (	read_data_1 	=> read_data_1,
        		read_data_2 	=> read_data_2,
        		Instruction 	=> Instruction,
				bubble_out		=> bubble_delay(0),--
        		read_data 		=> read_data,
				ALU_result 		=> ALU_result,
				RegWrite 		=> RegWrite,
				MemtoReg 		=> MemtoReg,
				RegDst 			=> RegDst,
				Sign_extend 	=> Sign_extend,
				IsSpecialAddr   => IsSpecialAddr,
				IsTEST=>IsTEST,
				addrOfIO=>addrOfIO,

        		clock 			=> clock,  
				reset 			=> reset );


   CTL:   control
	PORT MAP ( 	Opcode 			=> Instruction( 31 DOWNTO 26 ),
				RegDst 			=> RegDst,
				ALUSrc 			=> ALUSrc,
				MemtoReg 		=> MemtoReg,
				RegWrite 		=> RegWrite,
				MemRead 		=> MemRead,
				MemWrite 		=> MemWrite,
				Branch 			=> Branch,
				ALUop 			=> ALUop,
				Jump 			=> Jump,
				ICommand		=>ICommand,
				SLWCommand      =>SLWCommand,
				IsSWCommand     =>IsSWCommand,
				IsICommand  	=>IsICommand,
				clock 			=> clock,
				reset 			=> reset );

   EXE:  Execute
   	PORT MAP (	Read_data_1 	=> read_data_1,
             	Read_data_2 	=> read_data_2,
				Sign_extend 	=> Sign_extend,
                Function_opcode	=> Instruction( 5 DOWNTO 0 ),
				ALUOp 			=> ALUop,
				ALUSrc 			=> ALUSrc,
				Zero 			=> Zero,
                ALU_Result		=> ALU_Result,
				Add_Result 		=> Add_Result,
				PC_plus_4		=> PC_plus_4,
				ICommand		=>ICommand,
				SLWCommand      =>SLWCommand,
				IsSWCommand     =>IsSWCommand,
				IsICommand  	=>IsICommand,
				shiftValue      =>Instruction( 10 DOWNTO 6),
                Clock			=> clock,
				Reset			=> reset );

   MEM:  dmemory
	PORT MAP (	read_data 		=> read_data,
				address 		=>address_tmp,-- ALU_Result (9 DOWNTO 2)&"00",--jump memory address by 4
				write_data 		=> read_data_2,
				MemRead 		=> MemRead, 
				Memwrite 		=> MemWrite, 
				SpecialAddr     => SpecialAddr,
				SpecialData     => sw_0_7,
				IsSpecialAddr   =>IsSpecialAddr,
				Seven_Seg       =>Seven_Seg,
				PORT_LEDG=>PORT_LEDG,
				PORT_LEDR=>PORT_LEDR,
				addrOfIO=>addrOfIO,
                clock 			=> clock,  
				reset 			=> reset );
				
				
--==========================Convert from binary to hex= write data -> seven_seg===========================				
BCD0: BCD
	PORT MAP (
		Binary 	=> Seven_Seg( 3 downto 0 ),
		En 		=> the_one,
		Hex_out => ssg0_out );
	BCD1: BCD
	PORT MAP (
		Binary 	=> Seven_Seg( 7 downto 4 ),
		En 		=> the_one,
		Hex_out => ssg1_out );
	
	BCD2: BCD
	PORT MAP (
		Binary 	=> Seven_Seg( 11 downto 8 ),
		En 		=> the_one,
		Hex_out => ssg2_out );		
	
	BCD3: BCD
	PORT MAP (
		Binary 	=> Seven_Seg( 15 downto 12 ),
		En 		=> the_one,
		Hex_out => ssg3_out );
--=============================seven_segment display with DFF============================
  seg_signal_reg0: Ndff
    GENERIC MAP ( N => 7 )
	PORT MAP (	d 			=> ssg0_out,
				clk			=> clock,
				rst			=> reset,
				q			=> seg_signal_0 ); --goes to Idecode & control too
				
  seg_signal_reg1: Ndff
    GENERIC MAP ( N => 7 )
	PORT MAP (	d 			=> ssg1_out,
				clk			=> clock,
				rst			=> reset,
				q			=> seg_signal_1 ); --goes to Idecode & control too
				
  seg_signal_reg2: Ndff
    GENERIC MAP ( N => 7 )
	PORT MAP (	d 			=> ssg2_out,
				clk			=> clock,
				rst			=> reset,
				q			=> seg_signal_2 ); --goes to Idecode & control too

  seg_signal_reg3: Ndff
    GENERIC MAP ( N => 7 )
	PORT MAP (	d 			=> ssg3_out,
				clk			=> clock,
				rst			=> reset,
				q			=> seg_signal_3 ); --goes to Idecode & control too

END structure;
