 LIBRARY IEEE;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;
USE ieee.std_logic_unsigned.all;
USE work.aux_package.all;

ENTITY top_tb IS
	CONSTANT m : INTEGER := 8;
END top_tb;

architecture top_Testbench OF top_tb IS
SIGNAL rst,ena,clk: STD_LOGIC;
	SIGNAL din: STD_LOGIC_VECTOR (m-1 DOWNTO 0);
	SIGNAL cond : INTEGER range 0 to 3;
	SIGNAL	detector :  std_logic;
	SIGNAL	XX:  std_logic_vector(m-1 downto 0);
	SIGNAL	YY:  std_logic_vector(m-1 downto 0);

BEGIN

	L0 : top PORT MAP(rst,ena,clk,din,cond,detector,XX,YY);
		tb_ena : process
			begin 
			ena<='1';
			
			wait;
        end process tb_ena;
		
	tb_cond : process
		begin
				cond<=0;
			wait;
			
	end process tb_cond;

        tb_clk : process
			begin 
			clk<='1';
			wait for 5 us;
			clk<='0';
			wait for 5 us;
        end process tb_clk;
		
		tb_rst : process
			begin 
			rst<='1';
			wait for 5 us;
			rst<='0';
			wait;
        end process tb_rst;
		
		
    tb_din : process
		begin
			din <= "00000001";
			wait for 20 us;
			din <= "00000010";
			wait for 10 us;
			din <= "00000011"; 
			wait for 10 us;
			din <= "00000100";
			wait for 10 us;
			din <= "00001000";
			wait ;
        end process tb_din;
		

  
END top_Testbench;
